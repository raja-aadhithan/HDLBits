module top_module (input a,b,output q );
assign q = a&b;
endmodule
